module Instruction_Memory(read_addr, Instr_out);
    input [31:0]read_addr;
    output [31:0]Instr_out;
    reg [31:0]mem1[84:0];
initial begin
    mem1[0]  <= 32'b00000000000000001000001110110011; // add x7 , x1 , x0    
    mem1[4]  <= 32'b00000000000001010000000010110011; // add x1 , x10 , x0   
    mem1[8]  <= 32'b00000000000000111000010100110011; // add x10 , x7 , x0   
    mem1[12] <= 32'b00000000000000010000001110110011; // add x7 , x2 , x0  
    mem1[16] <= 32'b00000000000001011000000100110011; // add x2 , x11 , x0  
    mem1[20] <= 32'b00000000000000111000010110110011; // add x11 , x7 , x0
    mem1[24] <= 32'b00000000011101011000110000110011; // add x24 , x11 , x7
    mem1[28] <= 32'b00000001100011000000110000110011; // add x24 , x24, x24
    mem1[32] <= 32'b00000001010000000000101100010011; // addi x22 , x0 , 20
    mem1[36] <= 32'b00000000000000001010000100000011; // lw  x2,0(x1)
    mem1[40] <= 32'b00000000010100010000001000110011; // add x4 , x2 , x5
    mem1[44] <= 32'b00000000000000111000011010110011;
    mem1[48] <= 32'b00000001010000000000101100010011; //addi x22,x0,20
    mem1[52] <= 32'b00000001011011110010000000100011; //sw x22,0(x30)
    mem1[56] <= 32'b00000001000110000000001001100011; //beq x16,x17,4
    mem1[60] <= 32'b00000010100000000000101110010011; //addi x23,x0,40
    mem1[64] <= 32'b00000001100000000000110000010011; //addi x24,x0,24
    mem1[68] <= 32'b00000000000000001010001110000011; //lw x7,0(x5)
    mem1[72] <= 32'b00000001110011101111110010110011; //and x25, x29, x28
    mem1[76] <= 32'b00000001110011101101110110110011; //srl x27, x29, x28
    mem1[80] <= 32'b00000001110011101001111100110011; //sll x30, x29, x28
    mem1[84] <= 32'b00000000001011101001111110010011; //slli x31, x29, 2

end
assign Instr_out = mem1[read_addr];
endmodule