module ex_mem (
    input clk,
    input [2:0]wb,
    input [2:0]m,
    input [31:0]pc,
    input zero,
    input [31:0]alu_result,
    input [31:0]rs2,
    output [31:0]pc_out,
);
    
endmodule